module xor_gate_tb;

    reg A, B;
    wire Y;

    // Instantiate the XOR gate
    xor_gate uut (
        .A(A),
        .B(B),
        .Y(Y)
    );

    initial begin
        // Dump file for waveform
        $dumpfile("xor_gate.vcd");
        $dumpvars(0, xor_gate_tb);

        $display("A B | Y");
        $display("------");

        A = 0; B = 0; #10;
        A = 0; B = 1; #10;
        A = 1; B = 0; #10;
        A = 1; B = 1; #10;

        $finish;
    end

endmodule